library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity bancoRegistradores is
  port (
    HAB_ESCRITA_REG: in  std_logic;
    END1        : in  std_logic_vector(4 downto 0);
    END2        : in  std_logic_vector(4 downto 0);
    END3        : in  std_logic_vector(4 downto 0);
    DADO_W_REG3 : in  std_logic_vector(31 downto 0);
    DADO_R_REG1 : out std_logic_vector(31 downto 0);
    DADO_R_REG2 : out std_logic_vector(31 downto 0)
  );
end entity;

architecture bancoRegistradoresArch of bancoRegistradores is
  begin
    signal reset_reg : std_logic_vector (31 downto 0) :=  (others => '0');
    signal enable_write: std_logic_vector (31 downto 0 := (others => '0');
    signal out_reg0, out_reg1, out_reg2, out_reg3, out_reg4, out_reg5, out_reg6, out_reg7, out_reg8, out_reg9, out_reg10, out_reg11, out_reg12, out_reg13, out_reg14, out_reg15, out_reg16, 
           out_reg17, out_reg18, out_reg19, out_reg20, out_reg21, out_reg22, out_reg23, out_reg24, out_reg25, out_reg26, out_reg27, out_reg28, out_reg29, out_reg30, out_reg31 : std_logic_vector;

    REG0: entity work.registradorGenerico port map(DIN => dado_escrito_reg_3, DOUT => out_reg0, ENABLE => enable_write(0), CLK => clk, RST => reset_reg(0));
    REG1: entity work.registradorGenerico port map(DIN => dado_escrito_reg_3, DOUT => out_reg1, ENABLE => enable_write(1), CLK => clk, RST => reset_reg(1));
    REG2: entity work.registradorGenerico port map(DIN => dado_escrito_reg_3, DOUT => out_reg2, ENABLE => enable_write(2), CLK => clk, RST => reset_reg(2));
    REG3: entity work.registradorGenerico port map(DIN => dado_escrito_reg_3, DOUT => out_reg3, ENABLE => enable_write(3), CLK => clk, RST => reset_reg(3));
    REG4: entity work.registradorGenerico port map(DIN => dado_escrito_reg_3, DOUT => out_reg4, ENABLE => enable_write(4), CLK => clk, RST => reset_reg(4));
    REG5: entity work.registradorGenerico port map(DIN => dado_escrito_reg_3, DOUT => out_reg5, ENABLE => enable_write(5), CLK => clk, RST => reset_reg(5));
    REG6: entity work.registradorGenerico port map(DIN => dado_escrito_reg_3, DOUT => out_reg6, ENABLE => enable_write(6), CLK => clk, RST => reset_reg(6));
    REG7: entity work.registradorGenerico port map(DIN => dado_escrito_reg_3, DOUT => out_reg7, ENABLE => enable_write(7), CLK => clk, RST => reset_reg(7));
    REG8: entity work.registradorGenerico port map(DIN => dado_escrito_reg_3, DOUT => out_reg8, ENABLE => enable_write(8), CLK => clk, RST => reset_reg(8));
    REG9: entity work.registradorGenerico port map(DIN => dado_escrito_reg_3, DOUT => out_reg9, ENABLE => enable_write(9), CLK => clk, RST => reset_reg(9));
    REG10: entity work.registradorGenerico port map(DIN => dado_escrito_reg_3, DOUT => out_reg10, ENABLE => enable_write(10), CLK => clk, RST => reset_reg(10));
    REG11: entity work.registradorGenerico port map(DIN => dado_escrito_reg_3, DOUT => out_reg11, ENABLE => enable_write(11), CLK => clk, RST => reset_reg(11));
    REG12: entity work.registradorGenerico port map(DIN => dado_escrito_reg_3, DOUT => out_reg12, ENABLE => enable_write(12), CLK => clk, RST => reset_reg(12));
    REG13: entity work.registradorGenerico port map(DIN => dado_escrito_reg_3, DOUT => out_reg13, ENABLE => enable_write(13), CLK => clk, RST => reset_reg(13));
    REG14: entity work.registradorGenerico port map(DIN => dado_escrito_reg_3, DOUT => out_reg14, ENABLE => enable_write(14), CLK => clk, RST => reset_reg(14));
    REG15: entity work.registradorGenerico port map(DIN => dado_escrito_reg_3, DOUT => out_reg15, ENABLE => enable_write(15), CLK => clk, RST => reset_reg(15));
    REG16: entity work.registradorGenerico port map(DIN => dado_escrito_reg_3, DOUT => out_reg16, ENABLE => enable_write(16), CLK => clk, RST => reset_reg(16));
    REG17: entity work.registradorGenerico port map(DIN => dado_escrito_reg_3, DOUT => out_reg17, ENABLE => enable_write(17), CLK => clk, RST => reset_reg(17));
    REG18: entity work.registradorGenerico port map(DIN => dado_escrito_reg_3, DOUT => out_reg18, ENABLE => enable_write(18), CLK => clk, RST => reset_reg(18));
    REG19: entity work.registradorGenerico port map(DIN => dado_escrito_reg_3, DOUT => out_reg19, ENABLE => enable_write(19), CLK => clk, RST => reset_reg(19));
    REG20: entity work.registradorGenerico port map(DIN => dado_escrito_reg_3, DOUT => out_reg20, ENABLE => enable_write(20), CLK => clk, RST => reset_reg(20));
    REG21: entity work.registradorGenerico port map(DIN => dado_escrito_reg_3, DOUT => out_reg21, ENABLE => enable_write(21), CLK => clk, RST => reset_reg(21));
    REG22: entity work.registradorGenerico port map(DIN => dado_escrito_reg_3, DOUT => out_reg22, ENABLE => enable_write(22), CLK => clk, RST => reset_reg(22));
    REG23: entity work.registradorGenerico port map(DIN => dado_escrito_reg_3, DOUT => out_reg23, ENABLE => enable_write(23), CLK => clk, RST => reset_reg(23));
    REG24: entity work.registradorGenerico port map(DIN => dado_escrito_reg_3, DOUT => out_reg24, ENABLE => enable_write(24), CLK => clk, RST => reset_reg(24));
    REG25: entity work.registradorGenerico port map(DIN => dado_escrito_reg_3, DOUT => out_reg25, ENABLE => enable_write(25), CLK => clk, RST => reset_reg(25));
    REG26: entity work.registradorGenerico port map(DIN => dado_escrito_reg_3, DOUT => out_reg26, ENABLE => enable_write(26), CLK => clk, RST => reset_reg(26));
    REG27: entity work.registradorGenerico port map(DIN => dado_escrito_reg_3, DOUT => out_reg27, ENABLE => enable_write(27), CLK => clk, RST => reset_reg(27));
    REG28: entity work.registradorGenerico port map(DIN => dado_escrito_reg_3, DOUT => out_reg28, ENABLE => enable_write(28), CLK => clk, RST => reset_reg(28));
    REG29: entity work.registradorGenerico port map(DIN => dado_escrito_reg_3, DOUT => out_reg29, ENABLE => enable_write(29), CLK => clk, RST => reset_reg(29));
    REG30: entity work.registradorGenerico port map(DIN => dado_escrito_reg_3, DOUT => out_reg30, ENABLE => enable_write(30), CLK => clk, RST => reset_reg(30));
    REG31: entity work.registradorGenerico port map(DIN => dado_escrito_reg_3, DOUT => out_reg31, ENABLE => enable_write(31), CLK => clk, RST => reset_reg(31));



end architecture;
