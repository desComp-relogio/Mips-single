library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity bancoRegistradores is
  port (
    HAB_ESCRITA_REG : in  std_logic;
    CLK             : in  std_logic;
    END1            : in  std_logic_vector(4 downto 0);
    END2            : in  std_logic_vector(4 downto 0);
    END3            : in  std_logic_vector(4 downto 0);
    DADO_W_REG3     : in  std_logic_vector(31 downto 0);
    DADO_R_REG1     : out std_logic_vector(31 downto 0);
    DADO_R_REG2     : out std_logic_vector(31 downto 0)
  );
end entity;

architecture bancoRegistradoresArch of bancoRegistradores is
  signal end3_convert: integer := to_integer(unsigned(END3));
  signal dado_lido_1, dado_lido_2: std_logic_vector (31 downto 0) := (others => '0');
  signal reset_reg : std_logic_vector (31 downto 0) := (others => '0');
  signal enable_write: std_logic_vector (31 downto 0) := (others => '0');
  signal out_reg0, out_reg1, out_reg2, out_reg3, out_reg4, out_reg5, out_reg6, out_reg7, out_reg8, out_reg9, out_reg10, out_reg11, out_reg12, out_reg13, out_reg14, out_reg15, out_reg16, 
          out_reg17, out_reg18, out_reg19, out_reg20, out_reg21, out_reg22, out_reg23, out_reg24, out_reg25, out_reg26, out_reg27, out_reg28, out_reg29, out_reg30, out_reg31 : std_logic_vector(31 downto 0);

  begin
    REG0  : entity work.registradorGenerico port map(DIN => (others => '0'), DOUT => out_reg0, ENABLE => '1', CLK => CLK, RST => reset_reg(0));
    REG1  : entity work.registradorGenerico port map(DIN => DADO_W_REG3, DOUT => out_reg1, ENABLE => enable_write(1), CLK => CLK, RST => reset_reg(1));
    REG2  : entity work.registradorGenerico port map(DIN => DADO_W_REG3, DOUT => out_reg2, ENABLE => enable_write(2), CLK => CLK, RST => reset_reg(2));
    REG3  : entity work.registradorGenerico port map(DIN => DADO_W_REG3, DOUT => out_reg3, ENABLE => enable_write(3), CLK => CLK, RST => reset_reg(3));
    REG4  : entity work.registradorGenerico port map(DIN => DADO_W_REG3, DOUT => out_reg4, ENABLE => enable_write(4), CLK => CLK, RST => reset_reg(4));
    REG5  : entity work.registradorGenerico port map(DIN => DADO_W_REG3, DOUT => out_reg5, ENABLE => enable_write(5), CLK => CLK, RST => reset_reg(5));
    REG6  : entity work.registradorGenerico port map(DIN => DADO_W_REG3, DOUT => out_reg6, ENABLE => enable_write(6), CLK => CLK, RST => reset_reg(6));
    REG7  : entity work.registradorGenerico port map(DIN => DADO_W_REG3, DOUT => out_reg7, ENABLE => enable_write(7), CLK => CLK, RST => reset_reg(7));
    REG8  : entity work.registradorGenerico port map(DIN => DADO_W_REG3, DOUT => out_reg8, ENABLE => enable_write(8), CLK => CLK, RST => reset_reg(8));
    REG9  : entity work.registradorGenerico port map(DIN => DADO_W_REG3, DOUT => out_reg9, ENABLE => enable_write(9), CLK => CLK, RST => reset_reg(9));
    REG10 : entity work.registradorGenerico port map(DIN => DADO_W_REG3, DOUT => out_reg10, ENABLE => enable_write(10), CLK => CLK, RST => reset_reg(10));
    REG11 : entity work.registradorGenerico port map(DIN => DADO_W_REG3, DOUT => out_reg11, ENABLE => enable_write(11), CLK => CLK, RST => reset_reg(11));
    REG12 : entity work.registradorGenerico port map(DIN => DADO_W_REG3, DOUT => out_reg12, ENABLE => enable_write(12), CLK => CLK, RST => reset_reg(12));
    REG13 : entity work.registradorGenerico port map(DIN => DADO_W_REG3, DOUT => out_reg13, ENABLE => enable_write(13), CLK => CLK, RST => reset_reg(13));
    REG14 : entity work.registradorGenerico port map(DIN => DADO_W_REG3, DOUT => out_reg14, ENABLE => enable_write(14), CLK => CLK, RST => reset_reg(14));
    REG15 : entity work.registradorGenerico port map(DIN => DADO_W_REG3, DOUT => out_reg15, ENABLE => enable_write(15), CLK => CLK, RST => reset_reg(15));
    REG16 : entity work.registradorGenerico port map(DIN => DADO_W_REG3, DOUT => out_reg16, ENABLE => enable_write(16), CLK => CLK, RST => reset_reg(16));
    REG17 : entity work.registradorGenerico port map(DIN => DADO_W_REG3, DOUT => out_reg17, ENABLE => enable_write(17), CLK => CLK, RST => reset_reg(17));
    REG18 : entity work.registradorGenerico port map(DIN => DADO_W_REG3, DOUT => out_reg18, ENABLE => enable_write(18), CLK => CLK, RST => reset_reg(18));
    REG19 : entity work.registradorGenerico port map(DIN => DADO_W_REG3, DOUT => out_reg19, ENABLE => enable_write(19), CLK => CLK, RST => reset_reg(19));
    REG20 : entity work.registradorGenerico port map(DIN => DADO_W_REG3, DOUT => out_reg20, ENABLE => enable_write(20), CLK => CLK, RST => reset_reg(20));
    REG21 : entity work.registradorGenerico port map(DIN => DADO_W_REG3, DOUT => out_reg21, ENABLE => enable_write(21), CLK => CLK, RST => reset_reg(21));
    REG22 : entity work.registradorGenerico port map(DIN => DADO_W_REG3, DOUT => out_reg22, ENABLE => enable_write(22), CLK => CLK, RST => reset_reg(22));
    REG23 : entity work.registradorGenerico port map(DIN => DADO_W_REG3, DOUT => out_reg23, ENABLE => enable_write(23), CLK => CLK, RST => reset_reg(23));
    REG24 : entity work.registradorGenerico port map(DIN => DADO_W_REG3, DOUT => out_reg24, ENABLE => enable_write(24), CLK => CLK, RST => reset_reg(24));
    REG25 : entity work.registradorGenerico port map(DIN => DADO_W_REG3, DOUT => out_reg25, ENABLE => enable_write(25), CLK => CLK, RST => reset_reg(25));
    REG26 : entity work.registradorGenerico port map(DIN => DADO_W_REG3, DOUT => out_reg26, ENABLE => enable_write(26), CLK => CLK, RST => reset_reg(26));
    REG27 : entity work.registradorGenerico port map(DIN => DADO_W_REG3, DOUT => out_reg27, ENABLE => enable_write(27), CLK => CLK, RST => reset_reg(27));
    REG28 : entity work.registradorGenerico port map(DIN => DADO_W_REG3, DOUT => out_reg28, ENABLE => enable_write(28), CLK => CLK, RST => reset_reg(28));
    REG29 : entity work.registradorGenerico port map(DIN => DADO_W_REG3, DOUT => out_reg29, ENABLE => enable_write(29), CLK => CLK, RST => reset_reg(29));
    REG30 : entity work.registradorGenerico port map(DIN => DADO_W_REG3, DOUT => out_reg30, ENABLE => enable_write(30), CLK => CLK, RST => reset_reg(30));
    REG31 : entity work.registradorGenerico port map(DIN => DADO_W_REG3, DOUT => out_reg31, ENABLE => enable_write(31), CLK => CLK, RST => reset_reg(31));

    MUX_END_REG_1: entity work.mux32 port map(IN_0 => out_reg0, IN_1 => out_reg1, IN_2 => out_reg2, IN_3 => out_reg3, IN_4 => out_reg4, IN_5 => out_reg5, IN_6 => out_reg6, IN_7 => out_reg7, IN_8 => out_reg8, IN_9 => out_reg9, IN_10 => out_reg10, IN_11 => out_reg11, IN_12 => out_reg12, IN_13 => out_reg13, IN_14 => out_reg14, 
    IN_15 => out_reg15, IN_16 => out_reg16, IN_17 => out_reg17, IN_18 => out_reg18, IN_19 => out_reg19, IN_20 => out_reg20, IN_21 => out_reg21, IN_22 => out_reg22, IN_23 => out_reg23, IN_24 => out_reg24, IN_25 => out_reg25, IN_26 => out_reg26, IN_27 => out_reg27, IN_28 => out_reg28, IN_29 => out_reg29, IN_30 => out_reg30, IN_31 => out_reg31, SEL => END1, Q_OUT => dado_lido_1);
    DADO_R_REG1 <= dado_lido_1; 

    MUX_END_REG_2: entity work.mux32 port map(IN_0 => out_reg0, IN_1 => out_reg1, IN_2 => out_reg2, IN_3 => out_reg3, IN_4 => out_reg4, IN_5 => out_reg5, IN_6 => out_reg6, IN_7 => out_reg7, IN_8 => out_reg8, IN_9 => out_reg9, IN_10 => out_reg10, IN_11 => out_reg11, IN_12 => out_reg12, IN_13 => out_reg13, IN_14 => out_reg14, 
    IN_15 => out_reg15, IN_16 => out_reg16, IN_17 => out_reg17, IN_18 => out_reg18, IN_19 => out_reg19, IN_20 => out_reg20, IN_21 => out_reg21, IN_22 => out_reg22, IN_23 => out_reg23, IN_24 => out_reg24, IN_25 => out_reg25, IN_26 => out_reg26, IN_27 => out_reg27, IN_28 => out_reg28, IN_29 => out_reg29, IN_30 => out_reg30, IN_31 => out_reg31, SEL => END2, Q_OUT => dado_lido_2);
    DADO_R_REG2 <= dado_lido_2; 

    process(END3) 
    begin
      enable_write <= (others => '0');
      enable_write(end3_convert) <= HAB_ESCRITA_REG;
    end process;   

end architecture;
